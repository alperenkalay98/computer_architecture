module constant_value_generator2 #(parameter D=8'b00000000)(out);
	output [7:0] out;
	assign out = D;
endmodule
