module constant_value_generator #(parameter D=3'b000)(out);
	output [2:0] out;
	assign out = D;
endmodule
